../../../TheSDK_generators/verilog/f2_dsp_tapein6.v