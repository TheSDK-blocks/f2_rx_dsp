../../../TheSDK_generators/verilog/f2_rx_dsp.v