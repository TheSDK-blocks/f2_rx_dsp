../../../TheSDK_generators/verilog/tb_f2_rx_dsp.v