../../../TheSDK_generators/verilog/tb_f2_dsp_tapein6.v